//Instruction Decode Unit 

