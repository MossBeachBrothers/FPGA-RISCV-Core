//Register File 
