//Branch Unit 

