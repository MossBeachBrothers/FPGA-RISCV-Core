//Arithmetic Logic Unit

