//Control Unit 

