//Program Counter 
