//Instruction Fetch Unit 
